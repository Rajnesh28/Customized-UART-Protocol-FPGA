LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE IEEE.NUMERIC_STD.all;


ENTITY BaudRateGenerator is
	PORT(   CLOCK_50 	: IN STD_LOGIC; 
			  KEY 		: IN STD_LOGIC_VECTOR(3 downto 0);  
			  
			  ENABLE		: OUT STD_LOGIC);
	END BaudRateGenerator;

ARCHITECTURE RTL OF BaudRateGenerator IS

	SIGNAL COUNTER : INTEGER RANGE 0 TO 164;
	
BEGIN
PROCESS(KEY(3), CLOCK_50) 
BEGIN

IF (KEY(3) = '0') THEN
	COUNTER <= 0;
	
ELSIF (RISING_EDGE(CLOCK_50)) THEN

	COUNTER <= COUNTER + 1;

	IF (COUNTER = 162) THEN
		ENABLE <= '1';
		COUNTER <= 0;

	ELSE
		ENABLE <= '0';

	END IF;
	
END IF;

END PROCESS;
END;
