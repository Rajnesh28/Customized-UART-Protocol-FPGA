LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
 
LIBRARY WORK;
USE WORK.ALL;

ENTITY UART IS
	PORT(   CLOCK_50 	: IN STD_LOGIC; -- the fast clock for spinning wheel
			  KEY 		: IN STD_LOGIC_VECTOR(3 downto 0);  -- includes slow_clock and reset
			  
			  UART_RTX  : IN STD_LOGIC;
			  UART_RTS  : IN STD_LOGIC;
			  
			  
			  UART_TXD	: OUT STD_LOGIC;
			  UART_CTS	: OUT STD_LOGIC);
END UART;


ARCHITECTURE structural OF UART IS

COMPONENT TRANSMITTER is
	PORT(   CLOCK_50 	: IN STD_LOGIC; 
			  KEY 		: IN STD_LOGIC_VECTOR(3 downto 0);  
			  
			  UART_TXD	: OUT STD_LOGIC;
			  UART_CTS	: OUT STD_LOGIC);
END COMPONENT;

COMPONENT RECEIVER is
	PORT(   CLOCK_50 	: IN STD_LOGIC;
			  KEY 		: IN STD_LOGIC_VECTOR(3 downto 0);  
			  
			  UART_RTX  : IN STD_LOGIC;
			  UART_RTS  : IN STD_LOGIC);
end COMPONENT;


BEGIN

UART_T: TRANSMITTER PORT MAP (CLOCK_50 => CLOCK_50, KEY => KEY, UART_TXD => UART_TXD, UART_CTS => UART_CTS);

UART_R: RECEIVER PORT MAP (CLOCK_50 => CLOCK_50, KEY => KEY, UART_RTX => UART_RTX, UART_RTS => UART_RTS);

END;
