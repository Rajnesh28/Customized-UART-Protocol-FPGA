--Rajnesh Joshi & Devon Sandhu
--ENSC 350
--Lab Group 28

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY RECEIVER IS
	PORT(
			  CLOCK_50 : IN STD_LOGIC; --50Mhz
			  KEY 		: IN STD_LOGIC_VECTOR(3 downto 0);  
			  
			  UART_RXD  : IN STD_LOGIC;
			  
			  UART_CTS  : OUT STD_LOGIC;
			  LEDG 		: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			  LEDR 		: OUT STD_LOGIC_VECTOR(17 DOWNTO 0)

);		
end RECEIVER;

architecture rtl of RECEIVER is


COMPONENT Clock_Divider IS
PORT(CLOCK_50  : IN STD_LOGIC;
		KEY      : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		clk_out  : OUT STD_LOGIC);
END COMPONENT;
	
--States
type STATE IS (IDLE, WAITPERIODS, READ_DATA, DISPLAY_LCD, TRANSMIT_MESSAGE); 
SIGNAL CURRENT_STATE : STATE := IDLE; 

SIGNAL CLOCK : STD_LOGIC;
SIGNAL REDO_TRANSMIT : STD_LOGIC := '0';
SIGNAL PARITY_T		: STD_LOGIC := '0';
SIGNAL DATA_R		: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL PARITY_R		: STD_LOGIC := '1';



BEGIN
  
ClockDivider : CLOCK_DIVIDER PORT MAP (CLOCK_50 => CLOCK_50, KEY => KEY, CLK_OUT=>CLOCK);
  
NEXT_LOGIC : PROCESS(CLOCK, KEY(3))
VARIABLE CYCLES 		: INTEGER RANGE 0 TO 4000;
VARIABLE DATA_CYCLES : INTEGER RANGE 0 TO 3000;
VARIABLE INDEX 		: INTEGER RANGE 0 TO 20;
VARIABLE DATA_R		: STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN

IF (KEY(3) = '0') THEN
	LEDG(0) <= '1';
	CURRENT_STATE <= IDLE;

ELSIF (RISING_EDGE(CLOCK)) THEN

	CASE CURRENT_STATE IS 

	WHEN IDLE =>
		LEDG(2) <= UART_RXD;
		LEDG(0) <= '0';
		LEDG(1) <= '0';
		
		CYCLES := 0;
		DATA_CYCLES := 0;
		INDEX := 0;
		UART_CTS <= '1';
		
		IF (UART_RXD = '1') THEN
			UART_CTS <= '0';
			CURRENT_STATE <= WAITPERIODS;
		ELSE 
			CURRENT_STATE <= IDLE;
		END IF;
	
	WHEN WAITPERIODS => 
		IF (CYCLES = 1954) THEN	
			PARITY_R <= UART_RXD; --Register the first messageBit
			CURRENT_STATE <= READ_DATA;
		ELSE 
			CYCLES := CYCLES + 1;
			CURRENT_STATE <= WAITPERIODS;
		END IF;

	WHEN READ_DATA =>
	
		IF (DATA_CYCLES = 1303) THEN
			
			IF (INDEX < 8) THEN
				DATA_R(INDEX) := UART_RXD;
				INDEX := INDEX + 1;

				DATA_CYCLES := 0;
				CURRENT_STATE <= READ_DATA;
				
			ELSIF (INDEX = 8) THEN--STOP BIT WHICH IS TECHNICALLY A 1
				DATA_CYCLES := 0;
				CURRENT_STATE <= DISPLAY_LCD;
				
				
			END IF;
			
		ELSE
			DATA_CYCLES := DATA_CYCLES + 1;
			CURRENT_STATE <= TRANSMIT_MESSAGE;
		END IF;

			
--		WHEN VERIFY_PARITY =>
--			IF (DATA_R(INDEX) = '1') THEN
--				PARITY_R <= NOT PARITY_R;
--			ELSE
--				PARITY_R <= PARITY_R;
--			END IF;
--			
--			IF (INDEX < 7)THEN
--				INDEX := INDEX + 1;
--				CURRENT_STATE <= VERIFY_PARITY;
--			ELSIF (PARITY_R = PARITY_T) THEN
--				CURRENT_STATE <= DISPLAY_LCD;
--			ELSE
--				REDO_TRANSMIT <= '1';
--				CURRENT_STATE <= IDLE;
--			END IF;
--			
	WHEN DISPLAY_LCD =>
		CURRENT_STATE <= TRANSMIT_MESSAGE;
		
	WHEN TRANSMIT_MESSAGE =>
		
		LEDR(7 DOWNTO 0) <= DATA_R;
		LEDG(1) <= '1';
		CURRENT_STATE <= TRANSMIT_MESSAGE;
		
	
	END CASE;
		
		
END IF;
END PROCESS;

END;