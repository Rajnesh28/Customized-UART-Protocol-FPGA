LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
 
LIBRARY WORK;
USE WORK.ALL;

ENTITY UART IS
	PORT(   CLOCK_50 	: IN STD_LOGIC; -- the fast clock for spinning wheel
			  KEY 		: IN STD_LOGIC_VECTOR(3 downto 0);  -- includes slow_clock and reset
			  DATA		: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			  UART_CTS	: OUT STD_LOGIC
	);
END UART;


ARCHITECTURE structural OF UART IS

COMPONENT TRANSMITTER is
     port(
		  KEY		  : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  CLOCK_50 : IN STD_LOGIC;
		  
		  LEDG	  : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		  UART_CTS : OUT STD_LOGIC;
		  UART_TXD : OUT STD_LOGIC); 
end COMPONENT;

COMPONENT RECEIVER is
  port(
		  KEY		  : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		  CLOCK_50 : IN STD_LOGIC;
        UART_RTS : IN STD_LOGIC;
		  UART_RTX : IN STD_LOGIC;--
		  
		  LEDG	  : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		  DATA	  : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);					
end COMPONENT;

SIGNAL TXD : STD_LOGIC;

BEGIN

UART_T: TRANSMITTER port map(CLOCK_50 => CLOCK_50, KEY => KEY, UART_TXD => TXD);
UART_R: RECEIVER port map(CLOCK_50 => CLOCK_50, KEY => KEY, UART_RTX => TXD, DATA => DATA, UART_CTS => UART_CTS);

END;
